ARRAY: DBL : 100
     0      45.3407163942888
     1      41.4204388118444
     2      153.315110669152
     3      767.065016444337
     4      61.731379973577
     5      519.303215909425
     6      929.149789702683
     7      220.515532987432
     8      204.562919775286
     9      88.9926632349345
    10      699.690989544471
    11      706.461273928388
    12      494.630914411801
    13      261.77851914511
    14      711.571271862635
    15      378.366195307284
    16      200.64452951804
    17      232.607609700694
    18      436.096239572436
    19      469.498493927297
    20      861.18743608761
    21      977.238324460219
    22      444.519202897567
    23      34.2430994074061
    24      523.771740274398
    25      31.6387917993771
    26      753.173772130708
    27      591.588200811105
    28      822.891032240768
    29      329.578870595237
    30      232.078094143457
    31      536.528269078829
    32      430.618407870931
    33      403.581086734115
    34      987.324740266113
    35      966.909652560442
    36      850.530583341853
    37      867.514226523933
    38      311.605187743718
    39      148.390408674437
    40      997.598591259494
    41      639.523298311757
    42      468.074725693127
    43      931.914724377876
    44      690.77261895443
    45      815.406767099819
    46      541.534646666392
    47      572.806522051248
    48      159.216115325324
    49      945.25027272536
    50      821.333695119868
    51      155.413879619638
    52      41.074767262244
    53      343.613376535295
    54      110.019428706737
    55      96.5382741282407
    56      518.773273340786
    57      22.4050385981822
    58      561.483719647622
    59      856.876117576322
    60      516.908105237832
    61      674.524732248171
    62      737.174895003985
    63      698.460331977559
    64      22.799546840973
    65      191.983756232999
    66      670.991008016742
    67      345.871737387903
    68      66.2902784842487
    69      140.710484767664
    70      921.117490120752
    71      221.656459486883
    72      380.114596048423
    73      586.015785851523
    74      167.312806550093
    75      26.3396874192821
    76      691.126455874707
    77      762.343886197705
    78      713.69532482405
    79      77.3243178042231
    80      589.809335577213
    81      925.503046217143
    82      929.697771523938
    83      430.446002832822
    84      505.969611232155
    85      831.255978826087
    86      919.236130043509
    87      601.637641248125
    88      723.836457228212
    89      519.336634557385
    90      490.817005974621
    91      161.419415455973
    92      976.115568529868
    93      574.360281496477
    94      273.251111280756
    95      531.427295660333
    96      698.558163223117
    97      667.049290922959
    98      97.4325421719963
    99      548.736284742475
ARRAY: DONE