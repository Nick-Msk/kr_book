ARRAY: INT : 100
     0	   616
     1	   371
     2	   224
     3	   233
     4	   653
     5	   165
     6	   744
     7	   159
     8	    47
     9	   661
    10	   124
    11	   949
    12	   484
    13	   621
    14	   914
    15	    17
    16	   593
    17	   721
    18	   496
    19	    53
    20	   441
    21	   519
    22	   771
    23	    65
    24	   442
    25	   977
    26	   467
    27	   329
    28	   445
    29	   743
    30	   205
    31	   171
    32	   372
    33	   939
    34	   964
    35	   254
    36	    70
    37	   123
    38	   526
    39	   160
    40	   517
    41	   105
    42	   841
    43	   368
    44	   423
    45	   327
    46	   713
    47	   576
    48	   871
    49	   758
    50	   836
    51	   699
    52	   389
    53	   935
    54	   605
    55	   362
    56	   539
    57	   455
    58	   401
    59	   240
    60	    83
    61	   421
    62	   472
    63	   289
    64	   104
    65	   216
    66	   802
    67	   527
    68	   668
    69	   863
    70	   243
    71	   711
    72	   263
    73	   382
    74	    81
    75	   459
    76	   232
    77	   795
    78	   491
    79	     3
    80	   266
    81	   664
    82	   425
    83	   186
    84	   963
    85	   134
    86	   795
    87	   946
    88	   171
    89	   606
    90	    63
    91	   347
    92	   292
    93	   509
    94	   825
    95	   834
    96	   726
    97	   329
    98	   802
    99	   631
ARRAY: DONE